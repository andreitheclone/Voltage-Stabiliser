** Profile: "SCHEMATIC1-test1"  [ c:\users\gutaa\desktop\p1_2024_434d_guta_andrei_petrisor_sers_n13_orcad\p1_2024_434d_guta_andrei_petrisor_sers_n13_pspice\schematics\proiect_cef2-pspicefiles\schematic1\test1.sim ] 

** Creating circuit file "test1.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
* Local Libraries :
* From [PSPICE NETLIST] section of C:\Users\gutaa\AppData\Roaming\SPB_Data\cdssetup\OrCAD_PSpice\17.2.0\PSpice.ini file:
.lib "nomd.lib" 

*Analysis directives: 
.DC LIN I_I1 0 0.9 0.01 
.OPTIONS ADVCONV
.PROBE64 V(alias(*)) I(alias(*)) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC "..\SCHEMATIC1.net" 


.END
